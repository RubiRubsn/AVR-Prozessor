LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package
-- ---------------------------------------------------------------------------------
PACKAGE pkg_instrmem IS

	TYPE t_instrMem IS ARRAY(0 TO 512 - 1) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	CONSTANT PROGMEM : t_instrMem := (
		"0000000000000000",
		"1110000011100001",
		"1110000011110000",
		"1110101000011011",
		"1000001100010000",
		"1110111100011111",
		"1000000100010000",
		"1110000000000001",
		"1110101000010001",
		"1110101100100001",
		"1001001100101111",
		"1001001100011111",
		"1001001100001111",
		"1001000100101111",
		"1001000100011111",
		"1001000100001111",

		OTHERS => (OTHERS => '0')
	);

END PACKAGE pkg_instrmem;
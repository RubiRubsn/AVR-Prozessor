LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package
-- ---------------------------------------------------------------------------------
PACKAGE pkg_instrmem IS

	TYPE t_instrMem IS ARRAY(0 TO 512 - 1) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	CONSTANT PROGMEM : t_instrMem := (
		"1100000001100110",
		"1001001111111111",
		"1001001111101111",
		"1110000011110000",
		"1110001111100101",
		"1000001001110000",
		"1110001111101000",
		"1000001001100000",
		"1001000111101111",
		"1001000111111111",
		"1001010100001000",
		"1001001111111111",
		"1001001111101111",
		"1110000011110000",
		"1110001111100011",
		"1000000000110000",
		"1110001111100110",
		"1000000001000000",
		"1001000111101111",
		"1001000111111111",
		"1001010100001000",
		"1001001110001111",
		"1001001110011111",
		"1001001110111111",
		"1001001110101111",
		"1001001111001111",
		"1110000011000000",
		"0010111110101100",
		"0010111110111100",
		"0010110110000011",
		"0010110110010100",
		"0011000010010000",
		"1111000001001001",
		"0011000010000000",
		"1111000000111001",
		"1001010110000110",
		"1111010000010000",
		"0000111110101001",
		"0001111110111100",
		"0000111110011001",
		"0001111111001100",
		"1100111111110111",
		"0010111001111011",
		"0010111001101010",
		"1001000111001111",
		"1001000110101111",
		"1001000110111111",
		"1001000110011111",
		"1001000110001111",
		"1001010100001000",
		"1101111111100010",
		"1101111111001101",
		"1100000000101100",
		"1100000000101011",
		"1100000000101010",
		"1001001100001111",
		"1001001100011111",
		"1110000000010000",
		"0010110100000011",
		"0000110100000100",
		"0001111100010001",
		"0010111001110001",
		"0010111001100000",
		"1101111111000001",
		"1001000100011111",
		"1001000100001111",
		"1100000000011110",
		"1100000000011101",
		"1001001111111111",
		"1001001111101111",
		"1001001100001111",
		"1001001101001111",
		"1001001100011111",
		"1110000011110000",
		"1110001111100000",
		"1000000100000000",
		"0001010100000101",
		"1111000010011001",
		"1110111100011111",
		"0010010100010101",
		"0010001100010000",
		"0010111001010000",
		"0010111101000001",
		"0111000001000001",
		"1111011101110001",
		"0010111101000001",
		"0111000101000000",
		"1111011011010001",
		"0010111101000001",
		"0111000001001000",
		"1111011011010001",
		"0010111101000001",
		"0111000001000100",
		"1111011011000001",
		"0010111101000001",
		"0111000001000010",
		"1111011010110001",
		"1001000100011111",
		"1001000101001111",
		"1001000100001111",
		"1001000111101111",
		"1001000111111111",
		"1001010100001000",
		"1110000000000000",
		"0010111001010000",
		"0010111001110000",
		"0010111001100000",
		"1101111110011111",
		"1101111111010111",
		"1100111111111101",

		OTHERS => (OTHERS => '0')
	);

END PACKAGE pkg_instrmem;
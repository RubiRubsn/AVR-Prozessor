LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package
-- ---------------------------------------------------------------------------------
PACKAGE pkg_instrmem IS

	TYPE t_instrMem IS ARRAY(0 TO 512 - 1) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	CONSTANT PROGMEM : t_instrMem := (
		"0000000000000000",
		"1110010011100001",
		"1110000011110000",
		"1110101000011011",
		"1110101100101010",
		"1110111100111111",
		"1001001100011111",
		"1001001100101111",
		"1001001100111111",
		"1001000100101111",
		"1001000100011111",
		"1001000100111111",
		"0000000000000000",

		OTHERS => (OTHERS => '0')
	);

END PACKAGE pkg_instrmem;
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package
-- ---------------------------------------------------------------------------------
PACKAGE pkg_instrmem IS

	TYPE t_instrMem IS ARRAY(0 TO 512 - 1) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	CONSTANT PROGMEM : t_instrMem := (
		"0000000000000000",
		"1110010011100001",
		"1110000011110000",
		"1110101000011011",
		"1000001100010000",
		"1110010011100010",
		"1110101100011010",
		"1000001100010000",
		"1110010011100011",
		"1110111100010000",
		"1000001100010000",
		"1110010011100100",
		"1110000100010001",
		"1000001100010000",
		"1110010011100000",
		"1110111100011111",
		"1000001100010000",
		"0000000000000000",

		OTHERS => (OTHERS => '0')
	);

END PACKAGE pkg_instrmem;
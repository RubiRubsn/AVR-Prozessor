LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package
-- ---------------------------------------------------------------------------------
PACKAGE pkg_instrmem IS

	TYPE t_instrMem IS ARRAY(0 TO 512 - 1) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	CONSTANT PROGMEM : t_instrMem := (
		"0000000000000000",
		"1110111100011111",
		"1110000000100100",
		"1110000000110011",
		"0010111000110001",
		"1110101000011011",
		"1110000100100010",
		"0101000100100000",
		"1110000100100010",
		"0110000100100010",
		"1110000100100010",
		"0111000100100000",

		OTHERS => (OTHERS => '0')
	);

END PACKAGE pkg_instrmem;
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- ---------------------------------------------------------------------------------
-- Memory initialisation package
-- ---------------------------------------------------------------------------------
PACKAGE pkg_instrmem IS

	TYPE t_instrMem IS ARRAY(0 TO 512 - 1) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	CONSTANT PROGMEM : t_instrMem := (
		"0000000000000000",
		"1110110100010101",
		"0010111000110001",
		"0000000000000000",
		"1110000100010001",
		"0000110100010011",
		"0000000000000000",
		"1110000100010001",
		"0000111100010001",
		"0000000000000000",
		"1110000100010001",
		"1001010100010011",
		"0000000000000000",
		"1110111100011111",
		"1110000000000011",
		"0000110100010011",
		"0001111100010000",
		"0000000000000000",
		"1110000100010001",
		"1110000000000011",
		"0000111100010000",
		"0001111100010001",
		"0000000000000000",
		"1110000100010001",
		"0001100100010011",
		"0000000000000000",
		"1110000100010001",
		"0001010100010011",
		"0000000000000000",
		"1110000100010001",
		"0010111100000001",
		"0001011100010000",
		"0000000000000000",
		"1110000100010001",
		"0101000100010000",
		"0000000000000000",
		"1110000100010001",
		"0011000100010001",
		"0000000000000000",
		"1110000100010001",
		"1001010100011010",
		"0000000000000000",
		"1110000100010001",
		"0010100100010011",
		"0000000000000000",
		"1110000100010001",
		"0110101000011011",
		"0000000000000000",
		"1110000100010001",
		"0010010100010011",
		"0000000000000000",
		"1110000100010001",
		"1001010100010000",
		"0000000000000000",
		"1110000100010001",
		"0010000100010011",
		"0000000000000000",
		"1110000100010001",
		"0111101000011011",
		"0000000000000000",
		"1110101000011011",
		"1001010100010101",
		"0000000000000000",
		"1110101000011011",
		"1001010100010110",
		"0000000000000000",

		OTHERS => (OTHERS => '0')
	);

END PACKAGE pkg_instrmem;